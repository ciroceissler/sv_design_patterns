interface class brake_behavior_interface;
  pure virtual function void brake();
endclass : brake_behavior_interface
