interface class ice_cream_interface;
  pure virtual function void functionallity();
endclass : ice_cream_interface
