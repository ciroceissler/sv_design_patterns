class func1;

  int value;

  function new(int value=15);
    this.value = value;
  endfunction : new

endclass : func1
