class func2;

  int value;

  function new(int value=11);
    this.value = value;
  endfunction : new

endclass : func2
